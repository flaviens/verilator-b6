module top(in_data, out_data
// ,signal000_
// ,signal001_
// ,signal002_
// ,signal003_
// ,signal004_
// ,signal005_
// ,signal006_
// ,signal007_
// ,signal008_
// ,signal009_
// ,signal010_
// ,signal011_
// ,signal012_
// ,signal013_
// ,signal014_
// ,signal015_
// ,signal016_
// ,signal017_
// ,signal018_
// ,signal019_
// ,signal020_
// ,signal021_
// ,signal022_
// ,signal023_
// ,signal024_
// ,signal025_
// ,signal026_
// ,signal027_
// ,signal028_
// ,signal029_
// ,signal030_
// ,signal031_
// ,signal032_
// ,signal033_
// ,signal034_
// ,signal035_
// ,signal036_
// ,signal037_
// ,signal038_
// ,signal039_
// ,signal040_
// ,signal041_
// ,signal042_
// ,signal043_
// ,signal044_
// ,signal045_
// ,signal046_
// ,signal047_
// ,signal048_
// ,signal049_
// ,signal050_
// ,signal051_
// ,signal052_
// ,signal053_
// ,signal054_
// ,signal055_
// ,signal056_
// ,signal057_
// ,signal058_
// ,signal059_
// ,signal060_
// ,signal061_
// ,signal062_
// ,signal063_
// ,signal064_
// ,signal065_
// ,signal066_
// ,signal067_
// ,signal068_
// ,signal069_
// ,signal070_
// ,signal071_
// ,signal072_
// ,signal073_
// ,signal074_
// ,signal075_
// ,signal076_
// ,signal077_
// ,signal078_
// ,signal079_
// ,signal080_
// ,signal081_
// ,signal082_
// ,signal083_
// ,signal084_
// ,signal085_
// ,signal086_
// ,signal087_
// ,signal088_
// ,signal089_
// ,signal090_
// ,signal091_
// ,signal092_
// ,signal093_
// ,signal094_
// ,signal095_
// ,signal096_
// ,signal097_
// ,signal098_
// ,signal099_
// ,signal100_
// ,signal101_
// ,signal102_
// ,signal103_
// ,signal104_
// ,signal105_
// ,signal106_
// ,signal107_
// ,signal108_
// ,signal109_
// ,signal110_
// ,signal111_
// ,signal112_
// ,signal113_
// ,signal114_
// ,signal115_
// ,signal116_
// ,signal117_
// ,signal118_
// ,signal119_
// ,signal120_
// ,signal121_
// ,signal122_
// ,signal123_
// ,signal124_
// ,signal125_
// ,signal126_
// ,signal127_
// ,signal128_
// ,signal129_
// ,signal130_
// ,signal131_
// ,signal132_
// ,signal133_
// ,signal134_
// ,signal135_
// ,signal136_
// ,signal137_
// ,signal138_
// ,signal139_
// ,signal140_
// ,signal141_
// ,signal142_
// ,signal143_
// ,signal144_
// ,signal145_
// ,signal146_
// ,signal147_
// ,signal148_
// ,signal149_
// ,signal150_
// ,signal151_
// ,signal152_
// ,signal153_
// ,signal154_
// ,signal155_
// ,signal156_
// ,signal157_
// ,signal158_
// ,signal159_
// ,signal160_
// ,signal161_
// ,signal162_
// ,signal163_
// ,signal164_
// ,signal165_
// ,signal166_
// ,signal167_
// ,signal168_
// ,signal169_
// ,signal170_
// ,signal171_
// ,signal172_
// ,signal173_
// ,signal174_
// ,signal175_
// ,signal176_
// ,signal177_
// ,signal178_
// ,signal179_
// ,signal180_
// ,signal181_
// ,signal182_
// ,signal183_
// ,signal184_
// ,signal185_
);
  // output signal000_;
  // output signal001_;
  // output signal002_;
  // output signal003_;
  // output signal004_;
  // output signal005_;
  // output signal006_;
  // output signal007_;
  // output signal008_;
  // output signal009_;
  // output signal010_;
  // output signal011_;
  // output signal012_;
  // output signal013_;
  // output signal014_;
  // output signal015_;
  // output signal016_;
  // output signal017_;
  // output signal018_;
  // output signal019_;
  // output signal020_;
  // output signal021_;
  // output signal022_;
  // output signal023_;
  // output signal024_;
  // output signal025_;
  // output signal026_;
  // output signal027_;
  // output signal028_;
  // output signal029_;
  // output signal030_;
  // output signal031_;
  // output signal032_;
  // output signal033_;
  // output signal034_;
  // output signal035_;
  // output signal036_;
  // output signal037_;
  // output signal038_;
  // output signal039_;
  // output signal040_;
  // output signal041_;
  // output signal042_;
  // output signal043_;
  // output signal044_;
  // output signal045_;
  // output signal046_;
  // output signal047_;
  // output signal048_;
  // output signal049_;
  // output signal050_;
  // output signal051_;
  // output signal052_;
  // output signal053_;
  // output signal054_;
  // output signal055_;
  // output signal056_;
  // output signal057_;
  // output signal058_;
  // output signal059_;
  // output signal060_;
  // output signal061_;
  // output signal062_;
  // output signal063_;
  // output signal064_;
  // output signal065_;
  // output signal066_;
  // output signal067_;
  // output signal068_;
  // output signal069_;
  // output signal070_;
  // output signal071_;
  // output [281:0] signal072_;
  // output [281:0] signal073_;
  // output [281:0] signal074_;
  // output [14:0] signal075_;
  // output [14:0] signal076_;
  // output [14:0] signal077_;
  // output [238:0] signal078_;
  // output [238:0] signal079_;
  // output [61:0] signal080_;
  // output [61:0] signal081_;
  // output [61:0] signal082_;
  // output [72:0] signal083_;
  // output [72:0] signal084_;
  // output [299:0] signal085_;
  // output [299:0] signal086_;
  // output [299:0] signal087_;
  // output [61:0] signal088_;
  // output [66:0] signal089_;
  // output [66:0] signal090_;
  // output [19:0] signal091_;
  // output [259:0] signal092_;
  // output [259:0] signal093_;
  // output [259:0] signal094_;
  // output [60:0] signal095_;
  // output [60:0] signal096_;
  // output [60:0] signal097_;
  // output [81:0] signal098_;
  // output [81:0] signal099_;
  // output [200:0] signal100_;
  // output [200:0] signal101_;
  // output [200:0] signal102_;
  // output [296:0] signal103_;
  // output [296:0] signal104_;
  // output [219:0] signal105_;
  // output [219:0] signal106_;
  // output [174:0] signal107_;
  // output [174:0] signal108_;
  // output [6:0] signal109_;
  // output [88:0] signal110_;
  // output signal111_;
  // output [21:0] signal112_;
  // output [50:0] signal113_;
  // output [50:0] signal114_;
  // output [4:0] signal115_;
  // output [4:0] signal116_;
  // output [205:0] signal117_;
  // output [205:0] signal118_;
  // output [223:0] signal119_;
  // output [223:0] signal120_;
  // output [52:0] signal121_;
  // output [13:0] signal122_;
  // output [13:0] signal123_;
  // output signal124_;
  // output [109:0] signal125_;
  // output [109:0] signal126_;
  // output [298:0] signal127_;
  // output [298:0] signal128_;
  // output signal129_;
  // output [229:0] signal130_;
  // output [229:0] signal131_;
  // output [29:0] signal132_;
  // output [176:0] signal133_;
  // output [193:0] signal134_;
  // output [223:0] signal135_;
  // output [223:0] signal136_;
  // output [130:0] signal137_;
  // output [144:0] signal138_;
  // output [77:0] signal139_;
  // output [259:0] signal140_;
  // output [299:0] signal141_;
  // output [299:0] signal142_;
  // output [275:0] signal143_;
  // output [225:0] signal144_;
  // output [63:0] signal145_;
  // output [29:0] signal146_;
  // output [289:0] signal147_;
  // output [83:0] signal148_;
  // output [271:0] signal149_;
  // output [187:0] signal150_;
  // output [282:0] signal151_;
  // output [282:0] signal152_;
  // output [282:0] signal153_;
  // output [180:0] signal154_;
  // output [271:0] signal155_;
  // output [78:0] signal156_;
  // output [240:0] signal157_;
  // output [142:0] signal158_;
  // output [124:0] signal159_;
  // output [273:0] signal160_;
  // output [273:0] signal161_;
  // output [224:0] signal162_;
  // output [224:0] signal163_;
  // output [262:0] signal164_;
  // output [262:0] signal165_;
  // output [35:0] signal166_;
  // output [274:0] signal167_;
  // output [171:0] signal168_;
  // output [201:0] signal169_;
  // output [289:0] signal170_;
  // output [82:0] signal171_;
  // output [247:0] signal172_;
  // output [86:0] signal173_;
  // output [152:0] signal174_;
  // output [247:0] signal175_;
  // output [36:0] signal176_;
  // output [295:0] signal177_;
  // output [235:0] signal178_;
  // output [214:0] signal179_;
  // output [146:0] signal180_;
  // output [157:0] signal181_;
  // output [144:0] signal182_;
  // output [206:0] signal183_;
  // output [218:0] signal184_;
  // output [291:0] signal185_;

  bit signal000_;
  bit signal001_;
  bit signal002_;
  bit signal003_;
  bit signal004_;
  bit signal005_;
  bit signal006_;
  bit signal007_;
  bit signal008_;
  bit signal009_;
  bit signal010_;
  bit signal011_;
  bit signal012_;
  bit signal013_;
  bit signal014_;
  bit signal015_;
  bit signal016_;
  bit signal017_;
  bit signal018_;
  bit signal019_;
  bit signal020_;
  bit signal021_;
  bit signal022_;
  bit signal023_;
  bit signal024_;
  bit signal025_;
  bit signal026_;
  bit signal027_;
  bit signal028_;
  bit signal029_;
  bit signal030_;
  bit signal031_;
  bit signal032_;
  bit signal033_;
  bit signal034_;
  bit signal035_;
  bit signal036_;
  bit signal037_;
  bit signal038_;
  bit signal039_;
  bit signal040_;
  bit signal041_;
  bit signal042_;
  bit signal043_;
  bit signal044_;
  bit signal045_;
  bit signal046_;
  bit signal047_;
  bit signal048_;
  bit signal049_;
  bit signal050_;
  bit signal051_;
  bit signal052_;
  bit signal053_;
  bit signal054_;
  bit signal055_;
  bit signal056_;
  bit signal057_;
  bit signal058_;
  bit signal059_;
  bit signal060_;
  bit signal061_;
  bit signal062_;
  bit signal063_;
  bit signal064_;
  bit signal065_;
  bit signal066_;
  bit signal067_;
  bit signal068_;
  bit signal069_;
  bit signal070_;
  bit signal071_;
  bit [281:0] signal072_;
  bit [281:0] signal073_;
  bit [281:0] signal074_;
  bit [14:0] signal075_;
  bit [14:0] signal076_;
  bit [14:0] signal077_;
  bit [238:0] signal078_;
  bit [238:0] signal079_;
  bit [61:0] signal080_;
  bit [61:0] signal081_;
  bit [61:0] signal082_;
  bit [72:0] signal083_;
  bit [72:0] signal084_;
  bit [299:0] signal085_;
  bit [299:0] signal086_;
  bit [299:0] signal087_;
  bit [61:0] signal088_;
  bit [66:0] signal089_;
  bit [66:0] signal090_;
  bit [19:0] signal091_;
  bit [259:0] signal092_;
  bit [259:0] signal093_;
  bit [259:0] signal094_;
  bit [60:0] signal095_;
  bit [60:0] signal096_;
  bit [60:0] signal097_;
  bit [81:0] signal098_;
  bit [81:0] signal099_;
  bit [200:0] signal100_;
  bit [200:0] signal101_;
  bit [200:0] signal102_;
  bit [296:0] signal103_;
  bit [296:0] signal104_;
  bit [219:0] signal105_;
  bit [219:0] signal106_;
  bit [174:0] signal107_;
  bit [174:0] signal108_;
  bit [6:0] signal109_;
  bit [88:0] signal110_;
  bit signal111_;
  bit [21:0] signal112_;
  bit [50:0] signal113_;
  bit [50:0] signal114_;
  bit [4:0] signal115_;
  bit [4:0] signal116_;
  bit [205:0] signal117_;
  bit [205:0] signal118_;
  bit [223:0] signal119_;
  bit [223:0] signal120_;
  bit [52:0] signal121_;
  bit [13:0] signal122_;
  bit [13:0] signal123_;
  bit signal124_;
  bit [109:0] signal125_;
  bit [109:0] signal126_;
  bit [298:0] signal127_;
  bit [298:0] signal128_;
  bit signal129_;
  bit [229:0] signal130_;
  bit [229:0] signal131_;
  bit [29:0] signal132_;
  bit [176:0] signal133_;
  bit [193:0] signal134_;
  bit [223:0] signal135_;
  bit [223:0] signal136_;
  bit [130:0] signal137_;
  bit [144:0] signal138_;
  bit [77:0] signal139_;
  bit [259:0] signal140_;
  bit [299:0] signal141_;
  bit [299:0] signal142_;
  bit [275:0] signal143_;
  bit [225:0] signal144_;
  bit [63:0] signal145_;
  bit [29:0] signal146_;
  bit [289:0] signal147_;
  bit [83:0] signal148_;
  bit [271:0] signal149_;
  bit [187:0] signal150_;
  bit [282:0] signal151_;
  bit [282:0] signal152_;
  bit [282:0] signal153_;
  bit [180:0] signal154_;
  bit [271:0] signal155_;
  bit [78:0] signal156_;
  bit [240:0] signal157_;
  bit [142:0] signal158_;
  bit [124:0] signal159_;
  bit [273:0] signal160_;
  bit [273:0] signal161_;
  bit [224:0] signal162_;
  bit [224:0] signal163_;
  bit [262:0] signal164_;
  bit [262:0] signal165_;
  bit [35:0] signal166_;
  bit [274:0] signal167_;
  bit [171:0] signal168_;
  bit [201:0] signal169_;
  bit [289:0] signal170_;
  bit [82:0] signal171_;
  bit [247:0] signal172_;
  bit [86:0] signal173_;
  bit [152:0] signal174_;
  bit [247:0] signal175_;
  bit [36:0] signal176_;
  bit [295:0] signal177_;
  bit [235:0] signal178_;
  bit [214:0] signal179_;
  bit [146:0] signal180_;
  bit [157:0] signal181_;
  bit [144:0] signal182_;
  bit [206:0] signal183_;
  bit [218:0] signal184_;
  bit [291:0] signal185_;
  input [287:0] in_data;
  bit [287:0] in_data;
  output [159:0] out_data;
  bit [159:0] out_data;
  assign signal000_ = ~signal001_;
  assign signal002_ = ~signal003_;
  assign signal006_ = ~((signal008_ | in_data[29]) & signal007_);
  assign signal009_ = ~((signal012_ | signal011_) & signal010_);
  assign signal021_ = ~((signal023_ | signal022_) & (in_data[231] | in_data[71]));
  assign signal027_ = ~((signal031_ | signal030_) & (signal029_ | signal028_));
  assign signal032_ = signal033_ | ~(signal008_);
  assign signal034_ = signal021_ | ~(signal033_);
  assign signal035_ = signal033_ | ~(signal036_);
  assign signal037_ = signal026_ | ~(signal000_);
  assign signal018_ = in_data[126] | ~(signal002_);
  assign signal042_ = signal022_ | signal023_;
  assign signal043_ = signal044_ | in_data[64];
  assign signal004_ = signal045_ | signal001_;
  assign signal017_ = signal047_ | signal046_;
  assign signal048_ = signal050_ ^ signal049_;
  assign signal051_ = signal001_ ^ signal004_;
  assign signal052_ = signal054_ ^ signal053_;
  assign signal056_ = signal058_ ^ signal057_;
  assign signal044_ = signal060_ ^ signal059_;
  assign signal063_ = ~(signal059_ ^ signal064_);
  assign signal058_ = ~(signal065_ ^ signal043_);
  assign signal038_ = ~(signal066_ ^ signal058_);
  assign signal067_ = ~(signal051_ ^ signal028_);
  assign signal068_ = ~(signal069_ ^ signal043_);
  assign signal072_ = { signal074_[281:155], signal051_, signal074_[153:131], signal057_, signal074_[129:83], signal060_, signal074_[81:0] } + signal073_;
  assign signal075_ = { signal077_[14:1], signal053_ } + signal076_;
  assign signal080_ = { signal082_[61:4], signal004_, signal059_, signal028_, signal001_ } & { signal081_[61:1], signal022_ };
  assign signal083_ = { signal084_[72:43], signal023_, signal084_[41:0] } & { signal074_[115:83], signal060_, signal074_[81:45], signal004_, signal021_ };
  assign signal085_ = { in_data[274:119], signal087_[143:142], signal073_[132:1], signal052_, signal034_, signal087_[7:3], signal026_, signal053_, signal087_[0] } & { signal086_[299:290], signal025_, signal086_[288:262], signal056_, signal033_, signal086_[259:217], signal069_, signal086_[215:126], signal012_, signal086_[124:0] };
  assign out_data[51:32] = signal086_[181:162] & { signal091_[19:5], signal087_[6], signal022_, signal091_[2], signal032_, signal021_ };
  assign { signal092_[259:201], signal074_[281:155], signal092_[73:0] } = { signal094_[259:195], signal073_[132:1], signal094_[62:61], signal014_, signal094_[59:1], signal004_ } / { 1'h1, signal080_[31:9], signal093_[235], signal051_, signal046_, signal051_, signal093_[231:154], signal030_, signal093_[152:149], signal093_[149], signal093_[231:154], signal030_, signal093_[152:150], signal001_, signal049_, signal051_, signal008_, signal080_ };
  assign { signal095_[60], signal019_, signal095_[58:0] } = { signal097_[60:4], signal020_, signal044_, signal009_, signal097_[0] } / { 1'h1, signal096_[59:1], signal028_ };
  assign { signal093_[231:154], signal030_, signal093_[152:150] } = { signal099_[81:71], signal010_, signal099_[69:65], signal082_[61:4], signal099_[6:2], signal021_, signal051_ } / { 1'h1, signal098_[80:0] };
  assign signal100_ = { signal102_[200:180], signal094_[259:195], signal102_[114:88], signal079_[238:162], signal102_[10:1], signal011_ } / { 1'h1, signal101_[199:132], signal073_[132:1] };
  assign signal087_[5] = { signal092_[256:201], signal074_[281:250], signal021_ } == { signal086_[17:7], signal059_, signal023_, signal110_[75], signal008_, signal028_, signal083_ };
  assign signal111_ = { signal093_[164:154], signal030_, signal052_, signal073_[0], signal106_[143], signal063_, signal112_[5:3], signal112_[5:3] } == signal079_[231:210];
  assign out_data[96] = { signal114_[50:21], signal071_, signal114_[19:6], signal087_[143], signal021_, signal048_, signal041_, signal010_, signal028_ } == { signal097_[41:4], signal113_[12:4], signal067_, signal015_, signal087_[143], signal053_ };
  assign signal093_[149] = { in_data[64:30], signal087_[3], signal059_, signal049_, signal010_, signal046_, signal000_, signal041_ } === { signal074_[144:131], signal057_, signal074_[129:105], signal023_, signal051_ };
  assign signal012_ = { signal074_[153:137], signal093_[231:154], signal030_, signal093_[152:150], signal080_, signal080_, signal120_[0] } === { signal119_[223:49], signal101_[199:151] };
  assign signal074_[0] = { signal103_[136:120], signal081_[61:40], signal051_, signal080_, signal004_, signal041_, signal083_, signal051_ } === { signal103_[218:120], signal093_[235], signal000_, signal083_, signal001_, signal087_[3], signal093_[235], signal120_[0] };
  assign signal073_[0] = { signal083_[57:6], signal121_[0] } === { signal079_[205:162], signal102_[10:4], signal017_, signal087_[6] };
  assign signal053_ = { signal123_[13:9], signal102_[200:195], signal023_, signal022_, signal051_ } === { signal122_[13:1], signal042_ };
  assign signal124_ = { signal126_[109:3], signal002_, signal126_[1], signal052_ } === { signal125_[109:90], signal087_[5], signal106_[143], signal080_, signal087_[5], signal110_[75], signal116_[1], signal059_, signal125_[21], signal006_, signal087_[7], signal075_, signal001_, signal010_, signal125_[1], signal073_[0] };
  assign signal129_ = { signal131_[229:1], signal027_ } === { signal130_[229:115], signal115_, signal130_[109:0] };
  assign signal011_ = in_data[187:158] >= { signal014_, signal094_[59:43], signal041_, signal028_, signal051_, signal093_[235], signal000_, signal132_[6], signal044_, signal028_, signal087_[3], signal044_, signal028_, signal008_ };
  assign signal125_[21] = { signal133_[176:128], signal073_[281:154] } >= { signal079_[115:103], signal108_[167:133], signal086_[299:290], signal025_, signal086_[288:262], signal108_[94:5], signal074_[0] };
  assign signal099_[69] = { signal134_[193:181], signal131_[229:55], signal001_, signal004_, signal004_, signal023_, signal132_[6], signal023_ } >= { signal084_[50:43], signal023_, signal084_[41:10], signal132_[6], signal074_[153:131], signal057_, signal074_[129:83], signal060_, signal074_[81:2] };
  assign signal040_ = { signal102_[195:180], signal094_[259:195], signal102_[114:88], signal079_[238:169], signal136_[45:33], signal047_, signal136_[31:2], signal087_[3], signal087_[4] } > { signal135_[223:5], signal052_, signal087_[4], signal051_, signal046_, signal125_[1] };
  assign signal106_[147] = { signal137_[130:69], signal021_, signal059_, signal137_[66], signal137_[66], signal137_[64], signal080_, signal093_[149], signal078_[95] } > { signal074_[248:155], signal092_[73:38], signal078_[95] };
  assign signal022_ = { signal139_[77:72], signal099_[81:78], signal099_[69:65], signal082_[61:4], signal099_[6:2] } > { signal094_[59:58], signal099_[69], signal059_, signal099_[68:65], signal082_[61:4], signal099_[6:2], signal033_, signal041_, signal000_, signal132_[6], signal049_, signal059_, signal051_ };
  assign out_data[0] = { signal118_[204:194], signal086_[124:0], signal048_, signal079_[0], signal099_[68:65], signal082_[61:4], signal099_[6:2], signal015_, signal104_[50:0], signal038_, signal021_, signal009_ } > { signal140_[259:218], signal078_[238:127], signal075_, signal140_[90:65], signal013_, signal140_[63:41], signal103_[237], signal129_, signal140_[38:6], signal005_, signal140_[4:0] };
  assign signal059_ = { signal142_[299:269], signal141_[299:276], signal142_[244:228], signal096_[59:1], signal142_[168:165], signal023_, signal028_, signal132_[6], signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1], signal023_ } <= { signal141_[299:276], signal000_, signal141_[274:264], signal134_[193:181], signal131_[229:1], signal141_[21:0] };
  assign signal028_ = { in_data[276:25], signal132_[6] } && { in_data[286:35], signal023_ };
  assign signal121_[0] = { signal086_[112:76], signal143_[238], signal051_, signal093_[149], signal006_, signal063_, signal132_[6], signal001_, signal118_[144:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1], signal093_[231:154], signal030_, signal093_[152:150], signal034_, signal021_, signal143_[238], signal011_, signal044_, signal143_[238] } && { signal131_[218:27], signal001_, signal093_[231:154], signal030_, signal093_[152:150], signal093_[235] };
  assign signal074_[1] = { signal118_[203:182], signal024_ } && signal106_[35:13];
  assign signal097_[0] = { signal122_[2], signal022_, signal001_, signal049_, signal003_, signal026_, signal087_[6], signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:150], signal088_[61:40], signal036_, signal088_[38:0], signal144_[87:54], signal104_[50:0], signal034_, signal087_[7], signal061_ } && { signal092_[256:201], signal074_[281:155], signal092_[73:32], signal087_[4] };
  assign signal061_ = ! { signal096_[50:14], signal093_[149], signal087_[3], signal006_, signal093_[235] };
  assign signal016_ = ! { signal119_[133:49], signal101_[199:136], signal028_, signal049_ };
  assign signal087_[4] = ! { signal142_[232:228], signal096_[59:52] };
  assign signal076_[0] = ! { signal131_[105:43], signal149_[208], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:31], signal118_[144:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1], signal021_, signal063_, signal145_[36], signal087_[142] };
  assign signal127_[137] = ! { signal093_[210:154], signal030_, signal093_[152:150], signal112_[5:3], signal051_, signal020_, signal106_[141], signal051_, signal086_[259:217], signal069_, signal086_[215:126], signal058_, signal016_, signal074_[0] };
  assign signal029_ = ! { signal150_[187:114], signal097_[60:4], signal113_[12:4], signal150_[47:5], signal116_[4], signal079_[161], signal132_[6], signal051_, signal003_ };
  assign signal132_[6] = { in_data[15:12], in_data, signal023_, signal023_ } || { signal128_[273:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:5], signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1], signal023_ };
  assign signal145_[31] = { signal131_[215:210], signal046_, signal074_[0], signal100_, signal093_[149], signal000_, signal001_, signal087_[3], signal033_, signal021_, signal051_, signal099_[68:65], signal082_[61:4], signal099_[6:2] } || { in_data[14:11], signal011_, signal151_[277:224], signal138_[144:85], signal098_[80:0], signal138_[3:1], signal151_[79:63], signal022_, signal074_[0], signal012_, signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:160], signal093_[149] };
  assign signal145_[0] = { signal092_[259:201], signal074_[281:270] } || { signal086_[115:47], signal028_, signal028_ };
  assign signal148_[13] = { signal042_, signal062_, signal035_, signal147_[0], signal046_, signal020_, signal104_[50:0], signal153_[225:223], signal133_[176:128], signal073_[281:133], signal153_[24:5], signal044_, signal127_[137], signal001_, signal021_, signal074_[0] } || { signal084_[24:0], signal128_[184:169], signal006_, signal038_, signal152_[239:166], signal125_[109:90], signal152_[145:0] };
  assign out_data[64] = { signal106_[110:62], signal076_[14:1], signal106_[47:37], signal154_[106:96], signal078_[94:0], signal012_ } || { signal104_[181:137], signal089_[66:47], signal073_[132:17] };
  assign signal015_ = { signal102_[189:180], signal094_[259:234], signal041_ } < { signal144_[194:187], signal139_[77:72], signal099_[81:71], signal144_[169:162], signal001_, signal054_, signal110_[75], signal073_[0] };
  assign signal087_[143] = { signal119_[210:49], signal101_[199:140] } < { signal118_[125:91], signal118_[204:182], signal024_, signal090_[66:57], signal010_, signal074_[153:131], signal057_, signal074_[129:83], signal060_, signal074_[81:2] };
  assign signal010_ = signal132_[6] & ~(signal028_);
  assign signal033_ = signal132_[6] & ~(signal001_);
  assign { signal155_[271:256], signal123_[13:9], signal102_[200:180], signal094_[259:195], signal102_[114:88], signal079_[238:162], signal102_[10:1], signal155_[50:0] } = { signal141_[272:264], signal134_[193:181], signal131_[229:1], signal141_[21:3], signal001_, signal044_ } % { 1'h1, in_data[274:90], signal093_[149], signal000_, signal093_[231:154], signal030_, signal093_[152:150], signal051_, signal000_ };
  assign { signal136_[45:33], signal047_, signal136_[31:2] } = { signal073_[174:133], signal120_[0], signal132_[6] } % { 1'h1, signal074_[138:131], signal057_, signal074_[129:96] };
  assign signal086_[124:0] = { signal138_[124:85], signal098_[80:0], signal138_[3:1], signal151_[79] } % { 1'h1, signal082_[50:31], signal021_, signal044_, signal159_[101], signal157_[240:216], signal064_, signal157_[214:182], signal159_[41:36], signal050_, signal159_[34:6], signal049_, signal010_, signal110_[75], signal023_, signal093_[235], signal117_[79] };
  assign { signal144_[159:150], signal088_[61:40], signal036_, signal088_[38:0], signal144_[87:54] } = { signal154_[106:101], signal159_[101], signal157_[240:216], signal064_, signal157_[214:182], signal159_[41:36], signal050_, signal159_[34:6], signal032_, signal008_, signal110_[75], signal021_ } * { signal092_[233:201], signal074_[281:213], signal042_, signal001_, signal116_[1], signal074_[0] };
  assign { signal160_[273:245], signal130_[229:115], signal115_, signal130_[109:0], signal160_[14:0] } = { signal072_[281:63], signal117_[79], signal048_, signal074_[1], signal015_, signal104_[50:0] } * { signal079_[78:64], signal028_, signal074_[0], signal037_, signal161_[255:254], signal119_[223:49], signal101_[199:132], signal161_[10:2], signal132_[6], signal132_[6] };
  assign signal073_[132:1] = signal051_ ? { signal151_[253:224], signal138_[144:85], signal098_[80:42], signal006_, signal044_, signal087_[3] } : { signal084_[37:0], signal128_[184:160], signal099_[68:65], signal082_[61:4], signal099_[6:2], signal006_, signal008_ };
  assign { signal164_[262:197], signal140_[259:218], signal078_[238:99], signal164_[14:0] } = signal126_[1] ? { signal094_[16:10], signal124_, signal165_[254:242], signal126_[109:3], signal165_[134:0] } : { signal151_[264:224], signal138_[144:128], signal106_[141], signal100_, signal066_, signal087_[142], signal049_ };
  assign signal062_ = { signal074_[227:155], signal092_[73:6], signal001_, signal145_[31] } != { signal126_[70:3], signal165_[134:60] };
  assign signal020_ = { signal155_[268:256], signal123_[13:9], signal102_[200:180], signal094_[259:195], signal102_[114:88], signal079_[238:162], signal102_[10:1], signal155_[50:28], signal112_[5:3], signal022_ } != { signal086_[106:28], signal145_[36], signal125_[1], signal056_, signal015_, signal111_, signal079_[160:1], signal042_ };
  assign signal093_[235] = { in_data[173:51], signal023_, signal074_[153:131], signal057_, signal074_[129:83], signal060_, signal074_[81:2], signal023_, signal001_ } != { signal084_[10:8], signal141_[274:264], signal134_[193:181], signal131_[229:1], signal141_[21:0] };
  assign signal137_[66] = { signal119_[87:56], signal073_[0], signal006_, signal010_, signal087_[142] } != { signal103_[256:238], signal156_[57:54], signal026_, signal166_[11], signal148_[13], signal026_, signal087_[0], signal148_[13], signal099_[69], signal108_[1], signal051_, signal021_, signal041_, signal105_[2], signal106_[143] };
  assign signal154_[106:96] = - signal094_[32:22];
  assign { signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1] } = - in_data[252:92];
  assign { signal141_[274:264], signal134_[193:181], signal131_[229:1], signal141_[21:0] } = - { signal141_[282:276], signal142_[244:228], signal096_[59:1], signal142_[168:165], signal167_[187:165], signal028_, signal028_, signal001_, signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1], signal028_ };
  assign signal054_ = { signal136_[36:33], signal047_, signal136_[31:17], signal010_ } !== { signal083_[66:48], signal120_[0], signal061_ };
  assign signal087_[7] = { signal142_[234:228], signal096_[59:23], signal086_[259:217], signal069_, signal086_[215:126], signal026_, signal087_[6], signal074_[1], signal043_, signal046_, signal159_[101], signal157_[240:216], signal064_, signal157_[214:182], signal159_[41:36], signal050_, signal159_[34:6], signal087_[3], signal075_ } !== { signal080_[45:39], in_data };
  assign signal049_ = { signal167_[170:165], signal168_[165:161], signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1] } !== { signal131_[193:23], signal001_ };
  assign signal087_[0] = { signal157_[221:216], signal064_, signal157_[214:207], signal099_[68:65], signal082_[61:4], signal099_[6:2], signal015_, signal117_[79], signal058_, signal035_, signal042_, signal100_, signal145_[0], signal051_, signal034_ } !== { signal151_[226:224], signal138_[144:134], signal028_, signal044_, signal160_[273:245], signal130_[229:115], signal115_, signal130_[109:0], signal160_[14:0], signal147_[0] };
  assign signal116_[4] = { signal152_[143:17], signal032_, signal062_, signal166_[11], signal016_, signal088_[48:40], signal036_, signal088_[38:0], signal144_[87:68], signal039_, signal087_[5] } !== { signal140_[36:16], signal169_[180:1], signal106_[147] };
  assign signal079_[160:1] = ~ { signal100_[190:35], signal006_, signal021_, signal032_, signal074_[0] };
  assign signal078_[94:0] = ~ { signal088_[19:0], signal144_[87:84], signal028_, signal076_[0], signal026_, signal099_[68:65], signal082_[61:4], signal099_[6:2], signal020_ };
  assign { signal106_[138:62], signal076_[14:1], signal106_[47:1] } = { signal079_[155:22], signal010_, signal011_, signal041_, signal016_ } | { signal119_[141:49], signal101_[199:161], signal044_, signal147_[0], signal006_, signal032_, signal028_, signal087_[3] };
  assign signal112_[5:3] = { signal049_, signal048_, signal048_ } ** { signal082_[42], signal116_[1], signal093_[149] };
  assign signal171_ = { signal157_[229:216], signal064_, signal157_[214:182], signal159_[41:36], signal050_, signal159_[34:7] } ** { signal125_[92:90], signal152_[145:66] };
  assign { signal172_[247:245], signal162_[224:99], signal031_, signal162_[97:35], signal172_[54:0] } = { signal165_[245:242], signal126_[109:3], signal165_[134:3], signal059_, signal021_, signal066_, signal001_, signal166_[11] } ** { signal072_[280:36], signal021_, signal099_[69], signal087_[5] };
  assign { signal108_[167:133], signal086_[299:290], signal025_, signal086_[288:262], signal108_[94:5] } = { signal074_[279:155], signal092_[73:36] } ** { signal151_[229:224], signal138_[144:85], signal098_[80:0], signal138_[3:1], signal151_[79:71], signal103_[237], signal137_[64], signal018_, signal002_ };
  assign signal143_[238] = & { signal103_[171:120], signal103_[58:53], signal081_[61:1] };
  assign signal026_ = & { signal117_[79], signal021_, signal131_[214], signal146_[29:25], signal146_[11:1], signal163_[77:61], signal163_[31:3], signal122_[13:1], signal121_[0], signal063_, signal043_, signal033_, signal032_, signal100_, signal001_ };
  assign signal103_[237] = & { signal017_, signal100_[100:32] };
  assign signal041_ = & { signal004_, signal099_[68:65], signal099_[6:2], signal082_[61:4], signal051_ };
  assign signal079_[161] = & { signal140_[90:65], signal140_[63:41], signal020_, signal019_, signal015_, signal013_, signal030_, signal040_, signal150_[47:5], signal126_[1], signal170_[62], signal097_[28:4], signal095_[60], signal095_[58:3], signal113_[12:4], signal056_, signal093_[231:154], signal093_[152:150] };
  assign signal008_ = | signal119_[161:67];
  assign signal137_[64] = | signal131_[194:43];
  assign signal108_[1] = | { signal104_[33:28], signal022_, signal103_[237], signal106_[141] };
  assign signal126_[1] = | { signal095_[47:23], signal044_, signal108_[167:133], signal086_[299:290], signal025_, signal086_[288:262], signal108_[94:5], signal041_ };
  assign signal003_ = | { signal118_[204:182], signal118_[144:91], signal117_[79], signal090_[66:48], signal090_[46:1], signal147_[0], signal024_, signal055_, signal073_[262:166], signal073_[0], signal121_[0] };
  assign signal039_ = | signal072_[97:10];
  assign signal120_[0] = ^ { signal174_[152:137], signal142_[299:269], signal141_[299:276], signal142_[244:228], signal080_, signal006_, signal093_[235], signal099_[69] };
  assign signal110_[75] = ^ { signal144_[212:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:78] };
  assign signal087_[6] = ^ { in_data[205:35], signal074_[0], signal011_, signal032_, signal054_, signal066_, signal028_, signal110_[75] };
  assign signal147_[0] = signal093_[235] & signal004_;
  assign signal106_[143] = signal034_ & signal100_[113];
  assign signal079_[0] = signal130_[28] & signal002_;
  assign { signal159_[101], signal157_[240:216], signal064_, signal157_[214:182], signal159_[41:36], signal050_, signal159_[34:6] } = { signal079_[219:162], signal102_[10:1], signal155_[50:25], signal021_, signal087_[3] } >> { signal103_[183:155], signal099_[68:65], signal082_[61:4], signal099_[6:2] };
  assign { signal175_[247:245], signal104_[296:274], signal070_, signal104_[272:137], signal089_[66:47], signal104_[116:52] } = { signal072_[244:1], signal145_[0], signal125_[1], signal004_, signal125_[21] } >> { signal073_[200:152], signal042_, signal086_[259:217], signal069_, signal086_[215:126], signal017_, signal166_[11], signal094_[62:61], signal014_, signal094_[59:1] };
  assign { signal176_[36:28], signal091_[19:5], signal176_[12:0] } = signal171_[54:18] >> { signal086_[61:39], signal154_[106:96], signal040_, signal108_[1], signal033_ };
  assign { signal103_[235:120], signal081_[61:1], signal103_[58:0] } = { signal178_[235:207], signal174_[152:137], signal142_[299:269], signal141_[299:276], signal142_[244:228], signal096_[59:5], signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:160], signal051_, signal051_, signal021_, signal044_, signal022_ } << { in_data[185:10], signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:160], signal022_ };
  assign { signal099_[68:65], signal082_[61:4], signal099_[6:2] } = { signal131_[126:61], signal044_ } << { signal084_[53:43], signal023_, signal084_[41:0], signal128_[184:183], signal028_, signal028_, signal028_, signal001_, signal044_, signal000_, signal049_, signal059_, signal051_, signal028_, signal059_ };
  assign { signal151_[277:224], signal138_[144:85], signal098_[80:0], signal138_[3:1], signal151_[79:63] } = { signal179_[214], signal178_[235:207], signal174_[152:137], signal142_[299:269], signal141_[299:276], signal142_[244:228], signal096_[59:1], signal142_[168:165], signal167_[187:165], signal168_[165:161], signal179_[5:3], signal051_, signal093_[235], signal001_ } >> { signal074_[142:131], signal057_, signal074_[129:83], signal060_, signal074_[81:9], signal044_, signal049_, signal099_[69], signal044_, signal028_, signal132_[6], signal000_, signal044_, signal028_, signal001_, signal049_, signal004_, signal051_, signal093_[235], signal099_[68:65], signal082_[61:4], signal099_[6:2] };
  assign { signal180_[146:142], signal109_[5:1], signal180_[136:96], signal108_[174:168], signal180_[88:0] } = { signal074_[262:155], signal092_[73:37], signal004_, signal008_ } >> { signal094_[238:195], signal102_[114:88], signal079_[238:166], signal044_, signal023_, signal137_[64] };
  assign { signal094_[62:61], signal014_, signal094_[59:1] } = { signal131_[39:1], signal141_[21:1], signal023_, signal049_ } >> { signal128_[282:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:36] };
  assign { signal181_[157:97], signal173_[86:1], signal181_[10:0] } = { signal094_[29:4], signal073_[132:1] } <<< signal100_[165:8];
  assign { signal182_[144:142], signal158_[141:135], signal103_[295:238], signal156_[57:1], signal158_[19:3], signal182_[2:0] } = { signal085_[169:154], signal058_, signal087_[6], signal086_[124:0], signal058_, signal127_[137] } <<< { signal107_[157:15], signal166_[11], signal087_[7] };
  assign { signal163_[77:61], signal146_[29:25], signal122_[13:1], signal146_[11:1], signal163_[31:3] } = { signal088_[40], signal036_, signal088_[38:0], signal144_[87:54] } >>> { signal181_[153:97], signal173_[86:69] };
  assign { signal170_[258:246], signal150_[187:114], signal097_[60:4], signal113_[12:4], signal150_[47:5], signal170_[62] } = { signal100_[200:9], signal042_, signal011_, signal120_[0], signal023_, signal026_ } >>> { signal090_[48], signal055_, signal090_[46:14], signal079_[160:1], signal066_, signal106_[143] };
  assign signal104_[50:0] = { signal098_[47:0], signal138_[3:1] } >>> { signal098_[72:26], signal008_, signal016_, signal023_, signal061_ };
  assign { signal183_[206:200], signal114_[50:21], signal071_, signal114_[19:6], signal183_[154:121], signal077_[14:1], signal183_[106:99], signal127_[298:224], signal183_[23:0] } = { signal134_[189:181], signal131_[229:32] } >>> { signal046_, signal118_[144:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1], signal094_[62:61], signal014_, signal094_[59:1] };
  assign { signal177_[248:242], signal135_[223:5], signal177_[22:0] } = { signal072_[226:38], signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:160], signal143_[238] } >>> { signal118_[114:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:26], signal145_[31], signal094_[62:61], signal014_, signal094_[59:1], signal159_[101], signal157_[240:216], signal064_, signal157_[214:182], signal159_[41:36], signal050_, signal159_[34:6], signal034_ };
  assign { signal140_[38:6], signal005_, signal140_[4:0] } = signal171_[73:35] >>> { signal100_[185:180], signal145_[29:1], signal026_, signal028_, signal037_, signal087_[5] };
  assign signal107_[157:0] = { signal160_[266:245], signal130_[229:226], signal093_[231:154], signal030_, signal093_[152:150], signal125_[1], signal136_[45:33], signal047_, signal136_[31:2], signal011_, signal087_[3], signal043_, signal001_, signal087_[142] } >>> { signal150_[163:114], signal097_[60:4], signal113_[12:4], signal150_[47:10], signal149_[208], signal087_[4], signal106_[143], signal106_[143] };
  assign { signal118_[144:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1] } = { signal092_[17:4], signal086_[124:0], signal110_[75], signal046_, signal093_[235], signal041_, signal044_ } - { signal180_[129:96], signal108_[174:173], signal143_[238], signal011_, signal046_, signal012_, signal016_, signal143_[238], signal087_[3], signal011_, signal051_, signal022_, signal147_[0], signal159_[101], signal157_[240:216], signal064_, signal157_[214:182], signal159_[41:36], signal050_, signal159_[34:6], signal008_ };
  assign signal169_[180:1] = { signal151_[266:224], signal138_[144:85], signal098_[80:78], signal083_, signal078_[95] } - { signal162_[210:99], signal031_, signal162_[97:35], signal172_[54:53], signal051_, signal137_[64] };
  assign { signal152_[239:166], signal125_[109:90], signal152_[145:0] } = { signal119_[221:49], signal101_[199:134], signal121_[0] } ~^ { signal161_[254], signal119_[223:49], signal101_[199:137], signal093_[149] };
  assign { signal074_[153:131], signal057_, signal074_[129:83], signal060_, signal074_[81:2] } = in_data[250:99] ~^ { in_data[211:62], signal028_, signal000_ };
  assign { signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:160] } = { signal074_[68:13], signal059_, signal028_, signal028_ } ~^ { signal084_[35:0], signal128_[184:163], signal044_ };
  assign { signal161_[255:254], signal119_[223:49], signal101_[199:132], signal161_[10:2] } = { signal074_[123:83], signal060_, signal074_[81:34], signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1], signal004_, signal051_, signal049_ } ^ { signal131_[219:139], signal001_, signal093_[235], signal004_, signal041_, signal033_, signal051_, signal000_, signal028_, signal041_, signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1], signal023_, signal051_, signal093_[235] };
  assign { signal184_[218:212], signal179_[214], signal178_[235:207], signal174_[152:137], signal142_[299:269], signal141_[299:276], signal142_[244:228], signal096_[59:1], signal142_[168:165], signal167_[187:165], signal168_[165:161], signal179_[5:3] } = { in_data[184:129], signal028_, signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1], signal023_ } ^ { in_data[230:14], signal023_, signal023_ };
  assign { signal153_[225:223], signal133_[176:128], signal073_[281:133], signal153_[24:5] } = { signal073_[88:27], signal181_[157:97], signal173_[86:1], signal181_[10:0], signal051_ } ^ { signal144_[198:193], signal151_[277:224], signal138_[144:85], signal098_[80:0], signal138_[3:1], signal151_[79:63] };
  assign { signal086_[259:217], signal069_, signal086_[215:126] } = { signal125_[91:90], signal152_[145:14] } ^ { signal118_[141:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:10], signal042_, signal000_ };
  assign { signal140_[90:65], signal013_, signal140_[63:41] } = { signal088_[13:0], signal144_[87:54], signal121_[0], signal137_[64] } ^ { signal074_[201:155], signal092_[73], signal110_[75], signal000_ };
  assign signal145_[29:1] = { signal118_[202:182], signal024_, signal090_[66], signal061_, signal120_[0], signal117_[79], signal026_, signal120_[0], signal043_ } ^ { signal181_[153:133], signal006_, signal099_[69], signal017_, signal028_, signal003_, signal058_, signal015_, signal010_ };
  assign { signal185_[291:139], signal137_[130:69], signal185_[76:0] } = { signal172_[245], signal162_[224:99], signal031_, signal162_[97:35], signal172_[54:39], signal171_, signal041_, signal051_ } ^ { signal079_[135:62], signal058_, signal093_[231:154], signal030_, signal093_[152:150], signal087_[0], signal073_[132:1], signal127_[137], signal087_[5] };
  assign { signal165_[254:242], signal126_[109:3], signal165_[134:0] } = { signal131_[177:1], signal141_[21:14], signal099_[68:65], signal082_[61:4], signal099_[6:2], signal004_, signal041_, signal132_[6] } ^ { in_data[273:22], signal132_[6], signal132_[6], signal044_ };
  assign signal001_ = ~((signal179_[5] & signal132_[6]) | in_data[57]);
  assign signal166_[11] = ~((signal180_[127] & signal006_) | signal094_[33]);
  assign signal046_ = ~((signal093_[235] & signal004_) | (signal011_ & signal051_));
  assign signal106_[141] = ~((signal051_ & signal087_[6]) | (signal155_[12] & signal093_[149]));
  assign signal091_[2] = ~((signal149_[208] & signal068_) | (signal093_[149] & signal170_[248]));
  assign signal117_[79] = signal041_ ? signal165_[49] : signal032_;
  assign signal066_ = signal028_ ? signal094_[25] : signal120_[0];
  assign signal145_[36] = signal048_ ? signal048_ : signal094_[61];
  assign signal149_[208] = signal061_ ? signal180_[130] : signal010_;
  assign signal125_[1] = signal092_[258] ? signal028_ : signal043_;
  assign signal105_[2] = signal087_[142] ? signal145_[36] : signal106_[91];
  assign signal087_[142] = ~(signal110_[75] & signal054_);
  assign signal087_[3] = ~(signal033_ & signal144_[207]);
  assign signal078_[95] = !(signal087_[5] ? signal041_ : signal074_[74]);
  assign signal116_[1] = ~(signal062_ | signal126_[51]);
  assign { signal074_[154], signal074_[130], signal074_[82] } = { signal051_, signal057_, signal060_ };
  assign signal077_[0] = signal053_;
  assign signal078_[98:96] = { signal063_, signal008_, signal044_ };
  assign signal081_[0] = signal022_;
  assign signal082_[3:0] = { signal004_, signal059_, signal028_, signal001_ };
  assign signal084_[42] = signal023_;
  assign { signal086_[289], signal086_[261:260], signal086_[216], signal086_[125] } = { signal025_, signal056_, signal033_, signal069_, signal012_ };
  assign { signal087_[299:144], signal087_[141:8], signal087_[2:1] } = { in_data[274:119], signal073_[132:1], signal052_, signal034_, signal026_, signal053_ };
  assign signal088_[39] = signal036_;
  assign signal089_[46:0] = signal073_[132:86];
  assign { signal090_[47], signal090_[0] } = { signal055_, signal021_ };
  assign { signal091_[4:3], signal091_[1:0] } = { signal087_[6], signal022_, signal032_, signal021_ };
  assign signal092_[200:74] = signal074_[281:155];
  assign { signal093_[259:236], signal093_[234:232], signal093_[153], signal093_[148:0] } = { 1'h1, signal080_[31:9], signal051_, signal046_, signal051_, signal030_, signal093_[149], signal093_[231:154], signal030_, signal093_[152:150], signal001_, signal049_, signal051_, signal008_, signal080_ };
  assign { signal094_[194:63], signal094_[60], signal094_[0] } = { signal073_[132:1], signal014_, signal004_ };
  assign signal095_[59] = signal019_;
  assign { signal096_[60], signal096_[0] } = { 1'h1, signal028_ };
  assign signal097_[3:1] = { signal020_, signal044_, signal009_ };
  assign signal098_[81] = 1'h1;
  assign { signal099_[70], signal099_[64:7], signal099_[1:0] } = { signal010_, signal082_[61:4], signal021_, signal051_ };
  assign { signal101_[200], signal101_[131:0] } = { 1'h1, signal073_[132:1] };
  assign { signal102_[179:115], signal102_[87:11], signal102_[0] } = { signal094_[259:195], signal079_[238:162], signal011_ };
  assign { signal103_[296], signal103_[236], signal103_[119:59] } = { 1'h1, signal091_[2], signal081_[61:1] };
  assign { signal104_[273], signal104_[136:117], signal104_[51] } = { signal070_, signal089_[66:47], signal020_ };
  assign { signal105_[219:3], signal105_[1:0] } = { 1'h1, signal103_[225:120], signal081_[61:1], signal103_[58:10], signal012_, signal046_ };
  assign { signal106_[219:148], signal106_[146], signal106_[144], signal106_[142], signal106_[140], signal106_[61:48], signal106_[0] } = { signal103_[226:155], signal009_, signal063_, signal035_, signal021_, signal076_[14:1], signal027_ };
  assign signal107_[174:158] = { 1'h1, signal100_[141:128], signal004_, signal087_[4] };
  assign { signal108_[132:95], signal108_[4], signal108_[2], signal108_[0] } = { signal086_[299:290], signal025_, signal086_[288:262], signal043_, signal010_, signal073_[0] };
  assign { signal109_[6], signal109_[0] } = { 1'h1, signal044_ };
  assign { signal110_[88:76], signal110_[74:0] } = { signal086_[17:7], signal059_, signal023_, signal008_, signal028_, signal083_ };
  assign { signal112_[21:6], signal112_[2:0] } = { signal093_[164:154], signal030_, signal052_, signal073_[0], signal106_[143], signal063_, signal112_[5:3] };
  assign { signal113_[50:13], signal113_[3:0] } = { signal097_[41:4], signal067_, signal015_, signal087_[143], signal053_ };
  assign { signal114_[20], signal114_[5:0] } = { signal071_, signal087_[143], signal021_, signal048_, signal041_, signal010_, signal028_ };
  assign { signal116_[3], signal116_[0] } = { signal046_, signal023_ };
  assign signal117_[85:80] = { signal003_, signal112_[5:3], signal010_, signal106_[145] };
  assign { signal118_[205], signal118_[181:145], signal118_[90:0] } = { signal063_, signal024_, signal090_[66:48], signal055_, signal090_[46:31], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1], signal021_ };
  assign signal119_[48:0] = signal101_[199:151];
  assign signal120_[223:1] = { signal074_[153:137], signal093_[231:154], signal030_, signal093_[152:150], signal080_, signal080_ };
  assign signal121_[52:1] = signal083_[57:6];
  assign signal122_[0] = signal042_;
  assign signal123_[8:0] = { signal102_[200:195], signal023_, signal022_, signal051_ };
  assign { signal125_[89:22], signal125_[20:2], signal125_[0] } = { signal087_[5], signal106_[143], signal080_, signal087_[5], signal110_[75], signal116_[1], signal059_, signal006_, signal087_[7], signal075_, signal001_, signal010_, signal073_[0] };
  assign { signal126_[2], signal126_[0] } = { signal002_, signal052_ };
  assign { signal127_[139:138], signal127_[136:1] } = { signal124_, signal106_[143], signal086_[259:217], signal069_, signal086_[215:126], signal087_[4], signal018_ };
  assign { signal128_[298], signal128_[279], signal128_[257:185], signal128_[149:148], signal128_[146:0] } = { signal045_, signal007_, signal084_[72:43], signal023_, signal084_[41:0], signal087_[6], signal108_[1], signal051_, signal118_[144:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1], signal105_[2], signal126_[1] };
  assign signal130_[114:110] = signal115_;
  assign signal131_[0] = signal027_;
  assign { signal132_[29:7], signal132_[5:0] } = { signal014_, signal094_[59:43], signal041_, signal028_, signal051_, signal093_[235], signal000_, signal044_, signal028_, signal087_[3], signal044_, signal028_, signal008_ };
  assign signal133_[127:0] = signal073_[281:154];
  assign signal134_[180:0] = { signal131_[229:55], signal001_, signal004_, signal004_, signal023_, signal132_[6], signal023_ };
  assign signal135_[4:0] = { signal052_, signal087_[4], signal051_, signal046_, signal125_[1] };
  assign { signal136_[223:46], signal136_[32], signal136_[1:0] } = { signal102_[195:180], signal094_[259:195], signal102_[114:88], signal079_[238:169], signal047_, signal087_[3], signal087_[4] };
  assign { signal137_[68:67], signal137_[65], signal137_[63:0] } = { signal021_, signal059_, signal137_[66], signal080_, signal093_[149], signal078_[95] };
  assign { signal138_[84:4], signal138_[0] } = { signal098_[80:0], signal087_[142] };
  assign signal139_[71:0] = { signal099_[81:78], signal099_[69:65], signal082_[61:4], signal099_[6:2] };
  assign { signal140_[217:91], signal140_[64], signal140_[40:39], signal140_[5] } = { signal078_[238:127], signal075_, signal013_, signal103_[237], signal129_, signal005_ };
  assign { signal141_[275], signal141_[263:22] } = { signal000_, signal134_[193:181], signal131_[229:1] };
  assign { signal142_[268:245], signal142_[227:169], signal142_[164:13], signal142_[0] } = { signal141_[299:276], signal096_[59:1], signal023_, signal028_, signal132_[6], signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal023_ };
  assign { signal143_[275:239], signal143_[237:0] } = { signal086_[112:76], signal051_, signal093_[149], signal006_, signal063_, signal132_[6], signal001_, signal118_[144:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1], signal093_[231:154], signal030_, signal093_[152:150], signal034_, signal021_, signal143_[238], signal011_, signal044_, signal143_[238] };
  assign { signal144_[225:219], signal144_[203], signal144_[186:170], signal144_[149:88], signal144_[53:0] } = { signal122_[2], signal022_, signal001_, signal049_, signal003_, signal026_, signal087_[6], signal065_, signal139_[77:72], signal099_[81:71], signal088_[61:40], signal036_, signal088_[38:0], signal104_[50:0], signal034_, signal087_[7], signal061_ };
  assign { signal145_[63:40], signal145_[38:37], signal145_[35:32], signal145_[30] } = { signal088_[50:40], signal036_, signal088_[38:27], signal037_, signal042_, signal041_, signal062_, signal028_, signal125_[1], signal028_ };
  assign { signal146_[24:12], signal146_[0] } = { signal122_[13:1], signal076_[0] };
  assign signal147_[289:1] = { signal107_[69:46], signal027_, signal001_, signal127_[223], signal092_[259:201], signal074_[281:155], signal092_[73:0], signal132_[6], signal137_[64] };
  assign { signal148_[83:14], signal148_[11], signal148_[9:4], signal148_[2:0] } = { signal099_[66:65], signal082_[61:4], signal099_[6:2], signal108_[3], signal087_[7], signal066_, signal125_[21], signal087_[4], signal018_, signal063_, signal127_[223], signal039_, signal040_, signal103_[237], signal012_, signal040_, signal127_[223], signal020_ };
  assign { signal149_[271:209], signal149_[207:0] } = { signal131_[105:43], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:31], signal118_[144:91], signal118_[204:182], signal024_, signal090_[66:48], signal055_, signal090_[46:1], signal021_, signal063_, signal145_[36], signal087_[142] };
  assign { signal150_[113:48], signal150_[4:0] } = { signal097_[60:4], signal113_[12:4], signal116_[4], signal079_[161], signal132_[6], signal051_, signal003_ };
  assign { signal151_[282:278], signal151_[223:80], signal151_[62:0] } = { in_data[14:11], signal011_, signal138_[144:85], signal098_[80:0], signal138_[3:1], signal022_, signal074_[0], signal012_, signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:160], signal093_[149] };
  assign { signal152_[282:240], signal152_[165:146] } = { signal084_[24:0], signal128_[184:169], signal006_, signal038_, signal125_[109:90] };
  assign { signal153_[282:226], signal153_[222:25], signal153_[4:0] } = { signal042_, signal062_, signal035_, signal147_[0], signal046_, signal020_, signal104_[50:0], signal133_[176:128], signal073_[281:133], signal044_, signal127_[137], signal001_, signal021_, signal074_[0] };
  assign { signal154_[180:107], signal154_[95:0] } = { signal106_[110:62], signal076_[14:1], signal106_[47:37], signal078_[94:0], signal012_ };
  assign signal155_[255:51] = { signal123_[13:9], signal102_[200:180], signal094_[259:195], signal102_[114:88], signal079_[238:162], signal102_[10:1] };
  assign { signal156_[78:58], signal156_[0] } = { signal103_[258:238], signal002_ };
  assign { signal157_[215], signal157_[181:0] } = { signal064_, signal020_, signal093_[149], signal110_[75], signal015_, signal011_, signal088_[48:40], signal036_, signal088_[38:0], signal144_[87:68], signal039_, signal087_[5], signal074_[1], signal044_, signal104_[50:0], signal108_[1], signal140_[90:65], signal013_, signal140_[63:41], signal033_, signal001_ };
  assign { signal158_[142], signal158_[134:20], signal158_[2:1] } = { 1'h1, signal103_[295:238], signal156_[57:1], signal046_, signal056_ };
  assign { signal159_[124:102], signal159_[100:42], signal159_[35], signal159_[5:0] } = { 1'h1, signal082_[50:31], signal021_, signal044_, signal157_[240:216], signal064_, signal157_[214:182], signal050_, signal049_, signal010_, signal110_[75], signal023_, signal093_[235], signal117_[79] };
  assign signal160_[244:15] = { signal130_[229:115], signal115_, signal130_[109:0] };
  assign { signal161_[273:256], signal161_[253:11], signal161_[1:0] } = { signal079_[78:64], signal028_, signal074_[0], signal037_, signal119_[223:49], signal101_[199:132], signal132_[6], signal132_[6] };
  assign { signal162_[98], signal162_[34:2], signal162_[0] } = { signal031_, signal132_[6], signal126_[1], signal087_[7], signal145_[29:1], signal079_[0], signal105_[2] };
  assign { signal163_[224:78], signal163_[60:32], signal163_[2:0] } = { signal079_[159:13], signal146_[29:25], signal122_[13:1], signal146_[11:1], signal106_[141], signal132_[6], signal034_ };
  assign signal164_[196:15] = { signal140_[259:218], signal078_[238:99] };
  assign { signal165_[262:255], signal165_[241:135] } = { signal094_[16:10], signal124_, signal126_[109:3] };
  assign { signal166_[35:12], signal166_[10:0] } = { signal103_[256:238], signal156_[57:54], signal026_, signal148_[13], signal026_, signal087_[0], signal148_[13], signal099_[69], signal108_[1], signal051_, signal021_, signal041_, signal105_[2], signal106_[143] };
  assign { signal167_[274:188], signal167_[164:0] } = { signal141_[282:276], signal142_[244:228], signal096_[59:1], signal142_[168:165], signal028_, signal028_, signal001_, signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1], signal028_ };
  assign { signal168_[171:166], signal168_[160:0] } = { signal167_[170:165], signal045_, signal128_[297:280], signal007_, signal128_[278:258], signal084_[72:43], signal023_, signal084_[41:0], signal128_[184:150], signal142_[12:1] };
  assign { signal169_[201:181], signal169_[0] } = { signal140_[36:16], signal106_[147] };
  assign { signal170_[289:259], signal170_[245:63], signal170_[61:0] } = { signal085_[194:166], signal074_[1], signal058_, signal150_[187:114], signal097_[60:4], signal113_[12:4], signal150_[47:5], signal015_, signal095_[60], signal019_, signal095_[58:0] };
  assign signal172_[244:55] = { signal162_[224:99], signal031_, signal162_[97:35] };
  assign signal173_[0] = signal051_;
  assign signal174_[136:0] = { signal142_[299:269], signal141_[299:276], signal142_[244:228], signal080_, signal006_, signal093_[235], signal099_[69] };
  assign signal175_[244:0] = { signal104_[296:274], signal070_, signal104_[272:137], signal089_[66:47], signal104_[116:52] };
  assign signal176_[27:13] = signal091_[19:5];
  assign { signal177_[295:249], signal177_[241:23] } = { signal093_[204:158], signal135_[223:5] };
  assign signal178_[206:0] = { signal174_[152:137], signal142_[299:269], signal141_[299:276], signal142_[244:228], signal096_[59:5], signal144_[218:204], signal065_, signal144_[202:187], signal139_[77:72], signal099_[81:71], signal144_[169:160], signal051_, signal051_, signal021_, signal044_, signal022_ };
  assign { signal179_[213:6], signal179_[2:0] } = { signal178_[235:207], signal174_[152:137], signal142_[299:269], signal141_[299:276], signal142_[244:228], signal096_[59:1], signal142_[168:165], signal167_[187:165], signal168_[165:161], signal051_, signal093_[235], signal001_ };
  assign { signal180_[141:137], signal180_[95:89] } = { signal109_[5:1], signal108_[174:168] };
  assign signal181_[96:11] = signal173_[86:1];
  assign signal182_[141:3] = { signal158_[141:135], signal103_[295:238], signal156_[57:1], signal158_[19:3] };
  assign { signal183_[199:155], signal183_[120:107], signal183_[98:24] } = { signal114_[50:21], signal071_, signal114_[19:6], signal077_[14:1], signal127_[298:224] };
  assign signal184_[211:0] = { signal179_[214], signal178_[235:207], signal174_[152:137], signal142_[299:269], signal141_[299:276], signal142_[244:228], signal096_[59:1], signal142_[168:165], signal167_[187:165], signal168_[165:161], signal179_[5:3] };
  assign signal185_[138:77] = signal137_[130:69];
endmodule
